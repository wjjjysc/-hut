module seg7(
    input [3:0] q, // 二进制输入
    output reg [0:6] s //段码输出
);

// 个位数码管译码
always @* begin
    case(q)
        0: s = 7'b0000001; // 0
        1: s = 7'b1001111; // 1
        2: s = 7'b0010010; // 2
        3: s = 7'b0000110; // 3
        4: s = 7'b1001100; // 4
        5: s = 7'b0100100; // 5
        6: s = 7'b0100000; // 6
        7: s = 7'b0001111; // 7
        8: s = 7'b0000000; // 8
        9: s = 7'b0000100; // 9
        default: s = 7'b1111111; // 熄灭
    endcase
end


endmodule